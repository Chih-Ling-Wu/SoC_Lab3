`timescale 1ns / 1ps

module fir 
#(
    parameter pADDR_WIDTH = 12,
    parameter pDATA_WIDTH = 32,
    parameter Tape_Num    = 11
)
(
    output  wire                     awready,
    output  wire                     wready,
    input   wire                     awvalid,
    input   wire [(pADDR_WIDTH-1):0] awaddr,
    input   wire                     wvalid,
    input   wire [(pDATA_WIDTH-1):0] wdata,
    output  wire                     arready,
    input   wire                     rready,
    input   wire                     arvalid,
    input   wire [(pADDR_WIDTH-1):0] araddr,
    output  wire                     rvalid,
    output  wire [(pDATA_WIDTH-1):0] rdata,    
    input   wire                     ss_tvalid, 
    input   wire [(pDATA_WIDTH-1):0] ss_tdata, 
    input   wire                     ss_tlast, 
    output  wire                     ss_tready, 
    input   wire                     sm_tready, 
    output  wire                     sm_tvalid, 
    output  wire [(pDATA_WIDTH-1):0] sm_tdata, 
    output  wire                     sm_tlast, 
    
    // BRAM for tap RAM
    output  wire [3:0]               tap_WE,
    output  wire                     tap_EN,
    output  wire [(pDATA_WIDTH-1):0] tap_Di,
    output  wire [(pADDR_WIDTH-1):0] tap_A,
    input   wire [(pDATA_WIDTH-1):0] tap_Do,

    // BRAM for data RAM
    output  wire [3:0]               data_WE,
    output  wire                     data_EN,
    output  wire [(pDATA_WIDTH-1):0] data_Di,
    output  wire [(pADDR_WIDTH-1):0] data_A,
    input   wire [(pDATA_WIDTH-1):0] data_Do,

    input   wire                     axis_clk,
    input   wire                     axis_rst_n
);

    // Internal signals and registers
    reg [31:0] shift_reg [9:0]; // Shift register implemented with SRAM (11 DW)
    reg [31:0] tap_coeff [10:0]; // Tap coefficients implemented with SRAM (11 DW)
    reg [31:0] accum;
    reg [31:0] output_data;
    reg [4:0] tap_ptr;
    reg [31:0] data_count;
    wire tap_wr_enable;
    reg ap_start;

    // Internal AXI-Lite Control Registers
    reg [31:0] len_write_data;
    reg len_write_enable;
    reg [31:0] len_read_data;
    reg [31:0] ap_start_read_data;
    reg ap_start_write_enable;
    reg [31:0] ap_done_write_data;
    reg ap_done_write_enable;
    reg i;
    reg sm_tvalid_reg;

    // Address map constants
    localparam ADDR_AP_CTRL = 12'h00;
    localparam ADDR_DATA_LENGTH = 12'h10;
    localparam ADDR_TAP_PARAMS_START = 12'h20;
    localparam ADDR_TAP_PARAMS_END = 12'hFF;

    // Synthesizable reset logic
    always @(posedge axis_clk or negedge axis_rst_n) begin
        if (!axis_rst_n) begin
            // Reset your module's registers and state here
            for (i = 0; i < 11; i = i + 1) begin
                shift_reg[i] <= 0;
                tap_coeff[i] <= 0;
            end
            accum <= 0;
            output_data <= 0;
            tap_ptr <= 0;
            data_count <= 0;
            len_write_data <= 0;
            len_write_enable <= 0;
            len_read_data <= 0;
            ap_start_read_data <= 0;
            ap_start <= 0;
        end
    end

    // AXI-Lite Control Logic
    always @(posedge axis_clk or negedge axis_rst_n) begin
        if (!axis_rst_n) begin
            // Reset control signals
        end else begin
            // AXI-Lite address decoding
            case(awaddr)
                ADDR_AP_CTRL: begin
                    if (awvalid && !ap_start) begin
                        ap_start <= 1;
                        ap_done_write_enable <= 0;
                    end
                end
                ADDR_DATA_LENGTH: begin
                    if (awvalid) begin
                        len_write_data <= wdata;
                        len_write_enable <= 1;
                    end
                end
                ADDR_TAP_PARAMS_START: begin
                    if (awvalid) begin
                        // Write to tap coefficient BRAM
                        tap_WE <= awaddr[3:0];
                        tap_EN <= awvalid;
                        tap_Di <= wdata;
                        tap_A <= awaddr[(pADDR_WIDTH-1):2];
                    end
                end
                default: begin
                    len_write_enable <= 0;
                end
            endcase
        end
    end

    // Shift register implementation using SRAM
    always @(posedge axis_clk or posedge axis_rst_n) begin
        if (!axis_rst_n) begin
            // Reset shift register
            for (i = 0; i < 11; i = i + 1) begin
                shift_reg[i] <= 0;
            end
        end else if (ap_start) begin
            // Reset shift register on ap_start
            for (i = 0; i < 11; i = i + 1) begin
                shift_reg[i] <= 0;
            end
        end else if (ss_tvalid) begin
            // Shift in data when valid
            for (i = 10; i > 0; i = i - 1) begin
                shift_reg[i] <= shift_reg[i - 1];
            end
            shift_reg[0] <= ss_tdata;
        end
    end

    // FIR filtering logic
    always @(posedge axis_clk or posedge axis_rst_n) begin
        if (!axis_rst_n) begin
            // Reset FIR filter
            accum <= 0;
            output_data <= 0;
            tap_ptr <= 0;
            data_count <= 0;
        end else if (ap_start) begin
            // Reset FIR filter on ap_start
            accum <= 0;
            output_data <= 0;
            tap_ptr <= 0;
            data_count <= 0;
        end else if (ss_tvalid) begin
            // FIR filtering logic when data is valid
            // Shift in data when valid
            for (i = 10; i > 0; i = i - 1) begin
                shift_reg[i] <= shift_reg[i - 1];
            end
            shift_reg[0] <= ss_tdata;

            // Multiply and accumulate
            accum <= accum + (shift_reg[0] * tap_coeff[tap_ptr]);
            tap_ptr <= tap_ptr + 1;

            // Output valid data when tap pointer reaches Tape_Num
            if (tap_ptr == Tape_Num) begin
                output_data <= accum;
                accum <= 0;
                tap_ptr <= 0;
                data_count <= data_count + 1;
            end
        end
    end

    // AXI-Stream Output Logic
    reg [0:11] sm_tdata_reg;    // Register for sm_tdata signal
    reg sm_tlast_reg;           // Register for sm_tlast signal

    // AXI-Stream output logic
    always @(posedge axis_clk or negedge axis_rst_n) begin
        if (!axis_rst_n) begin
            // Reset AXI-Stream output signals and registers
            sm_tvalid_reg <= 0;
            sm_tdata_reg <= 0;
            sm_tlast_reg <= 0;
        end else if (ap_start) begin
            // Reset AXI-Stream output on ap_start
            sm_tvalid_reg <= 0;
            sm_tdata_reg <= 0;
            sm_tlast_reg <= 0;
        end else begin
            // Update output data register
            sm_tvalid_reg <= (data_count < len_read_data);
            sm_tdata_reg <= output_data;
            sm_tlast_reg <= (data_count == len_read_data - 1);
        end
    end

    // Drive the output signals with registered values
    assign sm_tvalid = sm_tvalid_reg;
    assign sm_tdata = sm_tdata_reg;
    assign sm_tlast = sm_tlast_reg;

    // Implement your AXI-Lite read logic for ap_start here
    always @(posedge axis_clk or negedge axis_rst_n) begin
        if (!axis_rst_n) begin
            // Reset AXI-Lite read logic for ap_start
            ap_start_read_data <= 0;
        end else begin
            if (ap_start_write_enable) begin
                ap_start_read_data <= ap_done_write_data;
            end
        end
    end
endmodule
